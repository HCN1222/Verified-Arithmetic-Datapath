.SUBCKT mux D0 D1 S Y vdd vss
*.PININFO D0:I D1:I S:I vdd:I vss:I Y:O
MM7 net19 S vdd vdd P_18 W=1.5u L=180.00n m=1
MM4 D1 net19 Y vdd P_18 W=1.5u L=180.00n m=1
MM3 D0 S Y vdd P_18 W=1.5u L=180.00n m=1
MM6 net19 S vss vss N_18 W=500.0n L=180.00n m=1
MM5 D1 S Y vss N_18 W=500.0n L=180.00n m=1
MM0 D0 net19 Y vss N_18 W=500.0n L=180.00n m=1
.ENDS

.SUBCKT inv vdd vin vout vss
*.PININFO vdd:I vin:I vss:I vout:O
MM1 vout vin vss vss N_18 W=500.0n L=180.00n m=1
MM0 vout vin vdd vdd P_18 W=1.5u L=180.00n m=1
.ENDS

.SUBCKT DFF1 CLK D Q VDD VSS
*.PININFO CLK:I D:I Q:O QB:O VDD:B VSS:B
MCLK_INV3_N net27 net11 VSS VSS N_18 W=500.0n L=180.00n
MD_INV2_N net0128 net0132 VSS VSS N_18 W=500.0n L=180.00n
MD_INV1_N net0132 D VSS VSS N_18 W=500.0n L=180.00n
MCLK_INV1_N net0136 CLK VSS VSS N_18 W=500.0n L=180.00n
MCLK_INV2_N net11 net0136 VSS VSS N_18 W=500.0n L=180.00n
MINV3_N net22 net9 VSS VSS N_18 W=500.0n L=180.00n
MINV1_N net9 net5 VSS VSS N_18 W=500.0n L=180.00n
MINV2_N Q net10 VSS VSS N_18 W=500.0n L=180.00n
MINV4_N QB Q VSS VSS N_18 W=500.0n L=180.00n
MCLK4_N net10 net27 QB VSS N_18 W=500.0n L=180.00n
MCLK3_N net9 net11 net10 VSS N_18 W=500.0n L=180.00n
MCLK1_N net0128 net27 net5 VSS N_18 W=500.0n L=180.00n
MCLK2_N net5 net11 net22 VSS N_18 W=500.0n L=180.00n
MCLK1_P net0128 net11 net5 VDD P_18 W=1.5u L=180.00n
MCLK_INV3_P net27 net11 VDD VDD P_18 W=1.5u L=180.00n
MD_INV2_P net0128 net0132 VDD VDD P_18 W=1.5u L=180.00n
MD_INV1_P net0132 D VDD VDD P_18 W=1.5u L=180.00n
MCLK_INV1_P net0136 CLK VDD VDD P_18 W=1.5u L=180.00n
MCLK_INV2_P net11 net0136 VDD VDD P_18 W=1.5u L=180.00n
MINV3_P net22 net9 VDD VDD P_18 W=1.5u L=180.00n
MINV1_P net9 net5 VDD VDD P_18 W=1.5u L=180.00n
MINV4_P QB Q VDD VDD P_18 W=1.5u L=180.00n
MINV2_P Q net10 VDD VDD P_18 W=1.5u L=180.00n
MCLK4_P net10 net11 QB VDD P_18 W=1.5u L=180.00n
MCLK3_P net9 net27 net10 VDD P_18 W=1.5u L=180.00n
MCLK2_P net5 net27 net22 VDD P_18 W=1.5u L=180.00n
.ENDS

.SUBCKT sub1 CLK r_clear_bar input max big_input pre VDD VSS
Xmux1 max input big_input max_temp VDD VSS / mux
Xmux2 pre max_temp r_clear_bar next_max VDD VSS / mux
XDFF CLK next_max max VDD VSS / DFF1
.ENDS

.SUBCKT sub2 CLK r_clear_bar input min big_input pre VDD VSS
Xmux1 input min big_input min_temp VDD VSS / mux
Xmux2 pre min_temp r_clear_bar next_min VDD VSS / mux
XDFF CLK next_min min VDD VSS / DFF1
.ENDS

.SUBCKT sub3 CLK r_clear_bar acc_result acc pre VDD VSS
Xmux pre acc_result r_clear_bar next_acc VDD VSS / mux
XDFF CLK next_acc acc VDD VSS / DFF1
.ENDS

.SUBCKT FA_MUX VDD VSS A B CIN COUT SUM
XINV1 VDD A N1 VSS / inv
XINV2 VDD N2 N3 VSS / inv
XMUX1 A N1 B N2 VDD VSS / mux
XMUX2 N2 N3 CIN SUM VDD VSS / mux
XMUX3 VSS A B N4 VDD VSS / mux
XMUX4 A VDD B N5 VDD VSS / mux
XMUX5 N4 N5 CIN COUT VDD VSS / mux
.ENDS

.SUBCKT ADDER4 VDD VSS A0 A1 A2 A3 B0 B1 B2 B3 CIN COUT S0 S1 S2 S3
XFA0 VDD VSS A0 B0 CIN COUT0 S0 / FA_MUX
XFA1 VDD VSS A1 B1 COUT0 COUT1 S1 / FA_MUX
XFA2 VDD VSS A2 B2 COUT1 COUT2 S2 / FA_MUX
XFA3 VDD VSS A3 B3 COUT2 COUT S3 / FA_MUX
.ENDS

.SUBCKT ADDER16 VDD VSS A0 A1 A2 A3 A4 A5 A6 A7 A8 A9 A10 A11 A12 A13 A14 A15 B0 B1 B2 B3 B4 B5 B6 B7 B8 B9 B10 B11 B12 B13 B14 B15 CIN COUT S0 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13 S14 S15
XAD40 VDD VSS A0 A1 A2 A3 B0 B1 B2 B3 CIN COUT0 S0 S1 S2 S3 / ADDER4
XAD41 VDD VSS A4 A5 A6 A7 B4 B5 B6 B7 COUT0 COUT1 S4 S5 S6 S7 / ADDER4
XAD42 VDD VSS A8 A9 A10 A11 B8 B9 B10 B11 COUT1 COUT2 S8 S9 S10 S11 / ADDER4
XAD43 VDD VSS A12 A13 A14 A15 B12 B13 B14 B15 COUT2 COUT S12 S13 S14 S15 / ADDER4
.ENDS

.SUBCKT TOP VDD VSS CLEAR CLK A0 A1 A2 A3 A4 A5 A6 A7 A8 A9 A10 A11 A12 A13 A14 A15 ACC0 ACC1 ACC2 ACC3 ACC4 ACC5 ACC6 ACC7 ACC8 ACC9 ACC10 ACC11 ACC12 ACC13 ACC14 ACC15 MAX0 MAX1 MAX2 MAX3 MAX4 MAX5 MAX6 MAX7 MAX8 MAX9 MAX10 MAX11 MAX12 MAX13 MAX14 MAX15 MIN0 MIN1 MIN2 MIN3 MIN4 MIN5 MIN6 MIN7 MIN8 MIN9 MIN10 MIN11 MIN12 MIN13 MIN14 MIN15
XFFCLEAR CLK CLEAR R_CLEAR VDD VSS / DFF1
XFFCLEARBAR VDD R_CLEAR R_CLEAR_BAR VSS / inv
XFF0 CLK A0 RIN0 VDD VSS / DFF1
XFF1 CLK A1 RIN1 VDD VSS / DFF1
XFF2 CLK A2 RIN2 VDD VSS / DFF1
XFF3 CLK A3 RIN3 VDD VSS / DFF1
XFF4 CLK A4 RIN4 VDD VSS / DFF1
XFF5 CLK A5 RIN5 VDD VSS / DFF1
XFF6 CLK A6 RIN6 VDD VSS / DFF1
XFF7 CLK A7 RIN7 VDD VSS / DFF1
XFF8 CLK A8 RIN8 VDD VSS / DFF1
XFF9 CLK A9 RIN9 VDD VSS / DFF1
XFF10 CLK A10 RIN10 VDD VSS / DFF1
XFF11 CLK A11 RIN11 VDD VSS / DFF1
XFF12 CLK A12 RIN12 VDD VSS / DFF1
XFF13 CLK A13 RIN13 VDD VSS / DFF1
XFF14 CLK A14 RIN14 VDD VSS / DFF1
XFF15 CLK A15 RIN15 VDD VSS / DFF1
XACCADDER VDD VSS ACC0 ACC1 ACC2 ACC3 ACC4 ACC5 ACC6 ACC7 ACC8 ACC9 ACC10 ACC11 ACC12 ACC13 ACC14 ACC15 RIN0 RIN1 RIN2 RIN3 RIN4 RIN5 RIN6 RIN7 RIN8 RIN9 RIN10 RIN11 RIN12 RIN13 RIN14 RIN15 VSS ACCCOUT ACCS0 ACCS1 ACCS2 ACCS3 ACCS4 ACCS5 ACCS6 ACCS7 ACCS8 ACCS9 ACCS10 ACCS11 ACCS12 ACCS13 ACCS14 ACCS15 / ADDER16
XSUB30 CLK R_CLEAR_BAR ACCS0 ACC0 VSS VDD VSS / sub3
XSUB31 CLK R_CLEAR_BAR ACCS1 ACC1 VSS VDD VSS / sub3
XSUB32 CLK R_CLEAR_BAR ACCS2 ACC2 VSS VDD VSS / sub3
XSUB33 CLK R_CLEAR_BAR ACCS3 ACC3 VSS VDD VSS / sub3
XSUB34 CLK R_CLEAR_BAR ACCS4 ACC4 VSS VDD VSS / sub3
XSUB35 CLK R_CLEAR_BAR ACCS5 ACC5 VSS VDD VSS / sub3
XSUB36 CLK R_CLEAR_BAR ACCS6 ACC6 VSS VDD VSS / sub3
XSUB37 CLK R_CLEAR_BAR ACCS7 ACC7 VSS VDD VSS / sub3
XSUB38 CLK R_CLEAR_BAR ACCS8 ACC8 VSS VDD VSS / sub3
XSUB39 CLK R_CLEAR_BAR ACCS9 ACC9 VSS VDD VSS / sub3
XSUB310 CLK R_CLEAR_BAR ACCS10 ACC10 VSS VDD VSS / sub3
XSUB311 CLK R_CLEAR_BAR ACCS11 ACC11 VSS VDD VSS / sub3
XSUB312 CLK R_CLEAR_BAR ACCS12 ACC12 VSS VDD VSS / sub3
XSUB313 CLK R_CLEAR_BAR ACCS13 ACC13 VSS VDD VSS / sub3
XSUB314 CLK R_CLEAR_BAR ACCS14 ACC14 VSS VDD VSS / sub3
XSUB315 CLK R_CLEAR_BAR ACCS15 ACC15 VSS VDD VSS / sub3
XINV0 VDD RIN0 RB0 VSS / inv
XINV1 VDD RIN1 RB1 VSS / inv
XINV2 VDD RIN2 RB2 VSS / inv
XINV3 VDD RIN3 RB3 VSS / inv
XINV4 VDD RIN4 RB4 VSS / inv
XINV5 VDD RIN5 RB5 VSS / inv
XINV6 VDD RIN6 RB6 VSS / inv
XINV7 VDD RIN7 RB7 VSS / inv
XINV8 VDD RIN8 RB8 VSS / inv
XINV9 VDD RIN9 RB9 VSS / inv
XINV10 VDD RIN10 RB10 VSS / inv
XINV11 VDD RIN11 RB11 VSS / inv
XINV12 VDD RIN12 RB12 VSS / inv
XINV13 VDD RIN13 RB13 VSS / inv
XINV14 VDD RIN14 RB14 VSS / inv
XINV15 VDD RIN15 RB15 VSS / inv
XMINADDER VDD VSS MIN0 MIN1 MIN2 MIN3 MIN4 MIN5 MIN6 MIN7 MIN8 MIN9 MIN10 MIN11 MIN12 MIN13 MIN14 MIN15 RB0 RB1 RB2 RB3 RB4 RB5 RB6 RB7 RB8 RB9 RB10 RB11 RB12 RB13 RB14 RB15 VDD MINCOUT MINS0 MINS1 MINS2 MINS3 MINS4 MINS5 MINS6 MINS7 MINS8 MINS9 MINS10 MINS11 MINS12 MINS13 MINS14 MINS15 / ADDER16
XSUB20 CLK R_CLEAR_BAR RIN0 MIN0 MINS15 VDD VDD VSS / sub2
XSUB21 CLK R_CLEAR_BAR RIN1 MIN1 MINS15 VDD VDD VSS / sub2
XSUB22 CLK R_CLEAR_BAR RIN2 MIN2 MINS15 VDD VDD VSS / sub2
XSUB23 CLK R_CLEAR_BAR RIN3 MIN3 MINS15 VDD VDD VSS / sub2
XSUB24 CLK R_CLEAR_BAR RIN4 MIN4 MINS15 VDD VDD VSS / sub2
XSUB25 CLK R_CLEAR_BAR RIN5 MIN5 MINS15 VDD VDD VSS / sub2
XSUB26 CLK R_CLEAR_BAR RIN6 MIN6 MINS15 VDD VDD VSS / sub2
XSUB27 CLK R_CLEAR_BAR RIN7 MIN7 MINS15 VDD VDD VSS / sub2
XSUB28 CLK R_CLEAR_BAR RIN8 MIN8 MINS15 VDD VDD VSS / sub2
XSUB29 CLK R_CLEAR_BAR RIN9 MIN9 MINS15 VDD VDD VSS / sub2
XSUB210 CLK R_CLEAR_BAR RIN10 MIN10 MINS15 VDD VDD VSS / sub2
XSUB211 CLK R_CLEAR_BAR RIN11 MIN11 MINS15 VDD VDD VSS / sub2
XSUB212 CLK R_CLEAR_BAR RIN12 MIN12 MINS15 VDD VDD VSS / sub2
XSUB213 CLK R_CLEAR_BAR RIN13 MIN13 MINS15 VDD VDD VSS / sub2
XSUB214 CLK R_CLEAR_BAR RIN14 MIN14 MINS15 VDD VDD VSS / sub2
XSUB215 CLK R_CLEAR_BAR RIN15 MIN15 MINS15 VSS VDD VSS / sub2
XINV16 VDD RIN0 RBA0 VSS / inv
XINV17 VDD RIN1 RBA1 VSS / inv
XINV18 VDD RIN2 RBA2 VSS / inv
XINV19 VDD RIN3 RBA3 VSS / inv
XINV20 VDD RIN4 RBA4 VSS / inv
XINV21 VDD RIN5 RBA5 VSS / inv
XINV22 VDD RIN6 RBA6 VSS / inv
XINV23 VDD RIN7 RBA7 VSS / inv
XINV24 VDD RIN8 RBA8 VSS / inv
XINV25 VDD RIN9 RBA9 VSS / inv
XINV26 VDD RIN10 RBA10 VSS / inv
XINV27 VDD RIN11 RBA11 VSS / inv
XINV28 VDD RIN12 RBA12 VSS / inv
XINV29 VDD RIN13 RBA13 VSS / inv
XINV30 VDD RIN14 RBA14 VSS / inv
XINV31 VDD RIN15 RBA15 VSS / inv
XMAXADDER VDD VSS MAX0 MAX1 MAX2 MAX3 MAX4 MAX5 MAX6 MAX7 MAX8 MAX9 MAX10 MAX11 MAX12 MAX13 MAX14 MAX15 RBA0 RBA1 RBA2 RBA3 RBA4 RBA5 RBA6 RBA7 RBA8 RBA9 RBA10 RBA11 RBA12 RBA13 RBA14 RBA15 VDD MAXCOUT MAXS0 MAXS1 MAXS2 MAXS3 MAXS4 MAXS5 MAXS6 MAXS7 MAXS8 MAXS9 MAXS10 MAXS11 MAXS12 MAXS13 MAXS14 MAXS15 / ADDER16
XSUB10 CLK R_CLEAR_BAR RIN0 MAX0 MAXS15 VSS VDD VSS / sub1
XSUB11 CLK R_CLEAR_BAR RIN1 MAX1 MAXS15 VSS VDD VSS / sub1
XSUB12 CLK R_CLEAR_BAR RIN2 MAX2 MAXS15 VSS VDD VSS / sub1
XSUB13 CLK R_CLEAR_BAR RIN3 MAX3 MAXS15 VSS VDD VSS / sub1
XSUB14 CLK R_CLEAR_BAR RIN4 MAX4 MAXS15 VSS VDD VSS / sub1
XSUB15 CLK R_CLEAR_BAR RIN5 MAX5 MAXS15 VSS VDD VSS / sub1
XSUB16 CLK R_CLEAR_BAR RIN6 MAX6 MAXS15 VSS VDD VSS / sub1
XSUB17 CLK R_CLEAR_BAR RIN7 MAX7 MAXS15 VSS VDD VSS / sub1
XSUB18 CLK R_CLEAR_BAR RIN8 MAX8 MAXS15 VSS VDD VSS / sub1
XSUB19 CLK R_CLEAR_BAR RIN9 MAX9 MAXS15 VSS VDD VSS / sub1
XSUB110 CLK R_CLEAR_BAR RIN10 MAX10 MAXS15 VSS VDD VSS / sub1
XSUB111 CLK R_CLEAR_BAR RIN11 MAX11 MAXS15 VSS VDD VSS / sub1
XSUB112 CLK R_CLEAR_BAR RIN12 MAX12 MAXS15 VSS VDD VSS / sub1
XSUB113 CLK R_CLEAR_BAR RIN13 MAX13 MAXS15 VSS VDD VSS / sub1
XSUB114 CLK R_CLEAR_BAR RIN14 MAX14 MAXS15 VSS VDD VSS / sub1
XSUB115 CLK R_CLEAR_BAR RIN15 MAX15 MAXS15 VDD VDD VSS / sub1
.ENDS






